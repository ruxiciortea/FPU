library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity normalization_unit is
    Port ( 
        clk: in std_logic;
        performed_operation: in std_logic;
        data_in: in std_logic_vector(31 downto 0);
        data_out: out std_logic_vector(31 downto 0)
    );
end normalization_unit;

architecture Behavioral of normalization_unit is

begin


end Behavioral;
